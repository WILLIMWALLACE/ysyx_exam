module ysyx_22040365_if(
  input		inst,
  input		clk,
  input		rst,
//  input		clr,
  output reg	inst,


);










endmodule
